module Addiererzelle (
    input [5:0] A,
    input [5:0] B,
    input C_IN,           // Carry In (Uebertragseingang)
    output reg[5:0] S,    // Summe
    output reg C_OUT      // Carry Out (Uebertragsausgang)
);
//something happens here
endmodule
